module Striking_pulse_generator (
    input wire CLK,
    input wire EN_work,
    input wire [3:0] sec_low,
    input wire [3:0] sec_high,
    input wire [3:0] min_low,
    input wire [3:0] min_high,
    input wire [3:0] hour_low,
    input wire [3:0] hour_high,
    output reg Chime
);

reg isChime;

// always @(posedge CLK or negedge EN_work) begin
always @(CLK) begin
    if (EN_work == 1'b0) begin
		// if(hour_low != 4'b0000 || hour_high != 4'b0000) begin // hour != 00 01 10 11
			if ((sec_low < 4'b0011 && sec_high == 4'b0000) && min_low == 4'b0000 && min_high == 4'b0000) begin
				// �����ĵ�λС�� 3����ĸ�λΪ 0���ҷ��ӵĵ�λ�͸�λ��Ϊ 0
				isChime <= 1'b1;  // ����isChime Ϊ 1
			end else begin
				isChime <= 1'b0;  // ����������������������� isChime Ϊ 0
			end
		//end else begin
		//	isChime <= 1'b0;
		//end
    end else begin
        isChime <= 1'b0;  // ��� EN_work ��Ϊ 0������ isChime Ϊ 0
    end
    
    //Chime <= isChime;  // �� isChime ��ֵ���� Chime ���
    Chime <= isChime;
end


endmodule